`timescale 1ns / 1ps

module four_to_one_demux_tb;

    reg S0, S1, S2, S3;
    wire I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15;
    four_to_one_demux DUT (
        .S0(S0),
        .S1(S1),
        .S2(S2),
        .S3(S3),
        .I0(I0),
        .I1(I1),
        .I2(I2),
        .I3(I3),
        .I4(I4),
        .I5(I5),
        .I6(I6),
        .I7(I7),
        .I8(I8),
        .I9(I9),
        .I10(I10),
        .I11(I11),
        .I12(I12),
        .I13(I13),
        .I14(I14),
        .I15(I15)
    );

    initial begin
        S0 = 0;
        S1 = 0;
        S2 = 0;
        S3 = 0;
        #20;

        S0 = 0;
        S1 = 0;
        S2 = 0;
        S3 = 1;
        #20;

        S0 = 0;
        S1 = 0;
        S2 = 1;
        S3 = 0;
        #20;

        S0 = 0;
        S1 = 0;
        S2 = 1;
        S3 = 1;
        #20;

        S0 = 0;
        S1 = 1;
        S2 = 0;
        S3 = 0;
        #20;

        S0 = 0;
        S1 = 1;
        S2 = 0;
        S3 = 1;
        #20;

        S0 = 0;
        S1 = 1;
        S2 = 1;
        S3 = 0;
        #20;

        S0 = 0;
        S1 = 1;
        S2 = 1;
        S3 = 1;
        #20;

        S0 = 1;
        S1 = 0;
        S2 = 0;
        S3 = 0;
        #20;

        S0 = 1;
        S1 = 0;
        S2 = 0;
        S3 = 1;
        #20;

        S0 = 1;
        S1 = 0;
        S2 = 1;
        S3 = 0;
        #20;

        S0 = 1;
        S1 = 0;
        S2 = 1;
        S3 = 1;
        #20;

        S0 = 1;
        S1 = 1;
        S2 = 0;
        S3 = 0;
        #20;

        S0 = 1;
        S1 = 1;
        S2 = 0;
        S3 = 1;
        #20;

        S0 = 1;
        S1 = 1;
        S2 = 1;
        S3 = 0;
        #20;

        S0 = 1;
        S1 = 1;
        S2 = 1;
        S3 = 1;
        #20;

        $finish;
    end

endmodule